﻿<?xml version="1.0" encoding="utf-8"?>
<ArrayOfVehiclesBase xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance" xmlns:xsd="http://www.w3.org/2001/XMLSchema">
  <VehiclesBase xsi:type="HybridCar">
    <Distance>453</Distance>
    <FuelConsumptionPerKm>18</FuelConsumptionPerKm>
    <CoefficientOfHybridity>3</CoefficientOfHybridity>
  </VehiclesBase>
  <VehiclesBase xsi:type="Car">
    <Distance>920</Distance>
    <FuelConsumptionPerKm>21</FuelConsumptionPerKm>
  </VehiclesBase>
  <VehiclesBase xsi:type="Helicopter">
    <Distance>7773</Distance>
    <FuelConsumptionPerKm>65</FuelConsumptionPerKm>
    <CargoWeight>715</CargoWeight>
  </VehiclesBase>
  <VehiclesBase xsi:type="Helicopter">
    <Distance>2294</Distance>
    <FuelConsumptionPerKm>43</FuelConsumptionPerKm>
    <CargoWeight>368</CargoWeight>
  </VehiclesBase>
  <VehiclesBase xsi:type="HybridCar">
    <Distance>335</Distance>
    <FuelConsumptionPerKm>11</FuelConsumptionPerKm>
    <CoefficientOfHybridity>9</CoefficientOfHybridity>
  </VehiclesBase>
</ArrayOfVehiclesBase>