﻿<?xml version="1.0" encoding="utf-8"?>
<ArrayOfVehiclesBase xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance" xmlns:xsd="http://www.w3.org/2001/XMLSchema">
  <VehiclesBase xsi:type="Helicopter">
    <Distance>2кк</Distance>
    <FuelConsumptionPerKm>20</FuelConsumptionPerKm>
    <CargoWeight>567</CargoWeight>
  </VehiclesBase>
  <VehiclesBase xsi:type="Car">
    <Distance>894</Distance>
    <FuelConsumptionPerKm>6</FuelConsumptionPerKm>
  </VehiclesBase>
  <VehiclesBase xsi:type="HybridCar">
    <Distance>785</Distance>
    <FuelConsumptionPerKm>15</FuelConsumptionPerKm>
    <CoefficientOfHybridity>8</CoefficientOfHybridity>
  </VehiclesBase>
  <VehiclesBase xsi:type="HybridCar">
    <Distance>319</Distance>
    <FuelConsumptionPerKm>21</FuelConsumptionPerKm>
    <CoefficientOfHybridity>6</CoefficientOfHybridity>
  </VehiclesBase>
  <VehiclesBase xsi:type="HybridCar">
    <Distance>834</Distance>
    <FuelConsumptionPerKm>27</FuelConsumptionPerKm>
    <CoefficientOfHybridity>2</CoefficientOfHybridity>
  </VehiclesBase>
  <VehiclesBase xsi:type="Helicopter">
    <Distance>4687</Distance>
    <FuelConsumptionPerKm>38</FuelConsumptionPerKm>
    <CargoWeight>851</CargoWeight>
  </VehiclesBase>
</ArrayOfVehiclesBase>